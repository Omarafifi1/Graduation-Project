module tw_factor_rom #(parameter addr_width = 3 , data_width = 64)(
  output [data_width-1:0] psi_1,psi_2,psi_3,psi_4,psi_5,psi_6,psi_7,psi_8,psi_9,psi_10,psi_11,psi_12,psi_13,psi_14,psi_15
);




assign psi_1=  32'h1da0;
assign psi_2=  32'h6c0;
assign psi_3=  32'h556;
assign psi_4=  32'h167c;
assign psi_5=  32'h94d;
assign psi_6=  32'h1bf2;
assign psi_7=  32'h13a9;
assign psi_8=  32'hd37;
assign psi_9=  32'h854;
assign psi_10= 32'h247;
assign psi_11= 32'h1321;
assign psi_12= 32'h4bd;
assign psi_13= 32'h1473;
assign psi_14= 32'h1ab0;
assign psi_15= 32'h15a7;


endmodule