module barret_reduction #(parameter data_size = 64 , parameter prime_number = 7681 ,
parameter no_of_bits_of_prime_no = $clog2(prime_number) , parameter factor_approximate_div = (2**(2*no_of_bits_of_prime_no)) / prime_number )
(
input [(data_size*2)-1:0] X ,
output reg signed [data_size-1 : 0] X_reduction
);


reg [data_size-1 : 0] q ;
reg [data_size-1 : 0] q_bar ;
reg [data_size-1 : 0] r , r_stage1,r_stage2,r_stage3 ,r_stage4 ;


always @(*) begin
if (X < prime_number) begin
	X_reduction = X ;
end
else begin
	q = X >> no_of_bits_of_prime_no ;
	q_bar = (q*factor_approximate_div) >> no_of_bits_of_prime_no ;
	r = X - (q_bar * prime_number) ;
	if (r >= prime_number) 
	r_stage1=r-prime_number;
	else 
	r_stage1=r;

	if (r_stage1>=prime_number) 
	r_stage2=r_stage1-prime_number;
	else 
	r_stage2=r_stage1;

	

	X_reduction=r_stage2;
end
end
endmodule