module barret_reduction #(
    parameter data_size = 64,
    parameter prime_number = 7681,
    parameter no_of_bits_of_prime_no = $clog2(prime_number),
    parameter factor_approximate_div = (2**(2*no_of_bits_of_prime_no)) / prime_number
)(
input   [(data_size*2)-1:0] X,
input   clk,rst_n,
output  signed  [data_size-1:0] X_reduction
);

// Pipeline registers
reg [data_size-1:0] q, q_bar;
reg [data_size-1:0] r, r_stage1;
reg [(data_size*2)-1:0]x_reg1 , x_reg2 , x_reg3;

always @(posedge clk , negedge rst_n) begin
	if(!rst_n)begin
		x_reg1<=0;
		x_reg2<=0;
	end
	else begin
		x_reg1<=X;
		x_reg2<=x_reg1;
	end
end

always @(posedge clk , negedge rst_n) begin
	if(!rst_n) begin
		r_stage1 <=0 ;
		q <=0 ;
		q_bar<=0;
		r<=0;
	end

	else begin
		// Pipeline Stage 1: Compute q and q_bar
		q <= X >> (no_of_bits_of_prime_no);
		q_bar <= (q * factor_approximate_div) >> (no_of_bits_of_prime_no);

		// Pipeline Stage 2: Compute initial remainder
		r <= x_reg2 - (q_bar * prime_number);

		// Pipeline Stage 3: 
		if (r >= prime_number)
			r_stage1 <= r - prime_number;
		else
			r_stage1 <= r;

	end
end
assign X_reduction=(r_stage1 >= prime_number)?r_stage1- prime_number:r_stage1;
endmodule
