module control_unit(
	input clk , rst_n,
	input start,
	output reg buffer_out_mux_selector_stage1 , buffer_in_mux_selector_stage1,
	output reg buffer_out_mux_selector_stage2 , buffer_in_mux_selector_stage2,
	output reg buffer_out_mux_selector_stage3 , buffer_in_mux_selector_stage3,
	output reg tw_factor_2nd_stage_mux_sel,
	output reg [1:0]tw_factor_3rd_stage_mux_sel,
	output reg buffer_enable,
	output done_tick
);

reg [4:0]counter ;

always @(posedge clk , negedge rst_n) begin
	if(!rst_n) begin
		counter<=0;	
	end
	else if(start)begin
		counter<=counter+1;
	end
end

always @(*) begin
	case (counter)
		5'd0, 5'd1, 5'd2, 5'd3:begin
			{buffer_out_mux_selector_stage1 , buffer_in_mux_selector_stage1}=2'bx1;
		end
		5'd4,5'd5,5'd6,5'd7,
		5'd12,5'd13,5'd14,5'd15,
		5'd20, 5'd21, 5'd22, 5'd23, 5'd24, 5'd25, 5'd26, 5'd27, 5'd28, 5'd29, 5'd30, 5'd31:begin
			{buffer_out_mux_selector_stage1 , buffer_in_mux_selector_stage1}=2'bxx;
		end

		5'd8 ,5'd9, 5'd10, 5'd11:begin
			{buffer_out_mux_selector_stage1 , buffer_in_mux_selector_stage1}=2'b10;
		end
		5'd16 ,5'd17 ,5'd18 ,5'd19:begin
			{buffer_out_mux_selector_stage1 , buffer_in_mux_selector_stage1}=2'b0x;
		end
	endcase


	case (counter)
		5'd8, 5'd9 :begin
			{buffer_out_mux_selector_stage2 , buffer_in_mux_selector_stage2}=2'bx1;
		end
		5'd0,5'd1,5'd2,5'd3,5'd4,5'd5,5'd6,5'd7,
		5'd10 ,5'd11 ,5'd12,5'd13,
		5'd18 ,5'd19 ,5'd20, 5'd21,
		5'd26, 5'd27, 5'd28, 5'd29, 5'd30, 5'd31:begin
			{buffer_out_mux_selector_stage2 , buffer_in_mux_selector_stage2}=2'bxx;
		end

		5'd14 ,5'd15 ,5'd22 ,5'd23:begin
			{buffer_out_mux_selector_stage2 , buffer_in_mux_selector_stage2}=2'b10;
		end
		5'd24 ,5'd25:begin
			{buffer_out_mux_selector_stage2 , buffer_in_mux_selector_stage2}=2'b0x;
		end
		5'd16 , 5'd17:begin
			{buffer_out_mux_selector_stage2 , buffer_in_mux_selector_stage2}=2'b01;
		end
	endcase

	case (counter)
		5'd14, 5'd16, 5'd24 :begin
			{buffer_out_mux_selector_stage3 , buffer_in_mux_selector_stage3}=2'bx1;
		end
		5'd0,5'd1,5'd2,5'd3,5'd4,5'd5,5'd6,5'd7,
		5'd8,5'd9,5'd10 ,5'd11 ,5'd12,5'd13 ,5'd15 ,5'd17 ,5'd18 ,5'd23 ,5'd25 ,5'd26 ,5'd31:begin
			{buffer_out_mux_selector_stage3 , buffer_in_mux_selector_stage3}=2'bxx;
		end

		5'd19 ,5'd21 ,5'd27 ,5'd29:begin
			{buffer_out_mux_selector_stage3 , buffer_in_mux_selector_stage3}=2'b10;
		end
		5'd20 ,5'd28 ,5'd30:begin
			{buffer_out_mux_selector_stage3 , buffer_in_mux_selector_stage3}=2'b0x;
		end
		5'd22:begin
			{buffer_out_mux_selector_stage3 , buffer_in_mux_selector_stage3}=2'b01;
		end
	endcase

	case (counter)
		5'd18 ,5'd19 ,5'd20 ,5'd21 ,5'd22 ,5'd23 ,5'd24 ,5'd25 ,5'd26 ,5'd27 ,5'd28 ,5'd29 ,5'd30 ,5'd31:begin
			tw_factor_2nd_stage_mux_sel=1'd1;
		end 
		default: tw_factor_2nd_stage_mux_sel=1'd0;
	endcase

	case (counter)
		5'd17, 5'd18, 5'd19, 5'd20, 5'd21, 5'd22: tw_factor_3rd_stage_mux_sel=2'd1;
		5'd23 ,5'd24 : tw_factor_3rd_stage_mux_sel=2'd2;
		5'd25 ,5'd26 ,5'd27 ,5'd28 ,5'd29 ,5'd30 ,5'd31: tw_factor_3rd_stage_mux_sel=2'd3;
		default: tw_factor_3rd_stage_mux_sel=2'd0;
	endcase

	case (counter)
		5'd12, 5'd13, 5'd14, 5'd15:begin
			buffer_enable=1'b0;
		end

		default:begin
			buffer_enable=1'b1;
		end		

	endcase
end
assign done_tick=(counter==5'd30);
endmodule